module mips_cpu_harvard_tb;
	timeunit 1ns / 10ps;

	parameter RAM_INIT_FILE = "";
	parameter TIMEOUT_CYCLES = 1000;
	parameter integer REF_OUT = 0;
	logic OUTPUT;
	logic clk;
	logic rst;
	logic clk_enable;
	logic active;
	logic[31:0] register_v0;
	logic[31:0] data_address;
	logic[31:0] instr_address;
	logic data_write;
	logic data_read;
	logic[31:0] data_writedata;
	logic[31:0] instr_readdata;
	logic[31:0] data_readdata;
	integer data_file;
	integer scan_file;
	mips_cpu_iMemory #(RAM_INIT_FILE) iMemory(instr_address,instr_readdata);
	mips_cpu_dMemory dMemory(clk,data_address,data_write,data_read,data_writedata,data_readdata);
	mips_cpu_harvard harvardCpu(clk,rst,active,register_v0,clk_enable,instr_address,instr_readdata,data_address,data_write,data_read,data_writedata,data_readdata);

	initial begin
		clk = 0;
		repeat(TIMEOUT_CYCLES) begin
			#10
			clk = !clk;
			#10
			clk = !clk;
		end

		$fatal(2,"CPU Timed Out, Infinite Loop",TIMEOUT_CYCLES);
	end

	initial begin
		rst <= 0;
		clk_enable <= 1;
		@(posedge clk);
		rst <= 1;
		@(posedge clk);
		#1
		assert(!(data_read || data_write));

		rst <= 0;
		@(posedge clk);
		assert(active==1);
		else $display("CPU signal active != 1 after reset");


		while(active) begin
		 @(posedge clk);
		 assert(!(data_read && data_write));
		 if(data_write) begin
		 	assert(instr_address != data_address);
		 end
		 //$display("Tick");
		 //$display("instr_address : %32h, instr_readdata : %32h data_address: %32h data_writedata: %32h data_readdata : %32h read: %1b write: %1b",instr_address,instr_readdata,data_address,data_writedata,data_readdata,data_read,data_write);
		end
		//$display("Register V0: ",register_v0);
		//$display("Finished Running");
		//scan_file = $fscanf(REF_FILE, "%d\n", OUTPUT);
		if(register_v0 != REF_OUT) begin
			$fatal(1,"Reference Outputs do not match Testbench Output: %h, %h", register_v0,REF_OUT);
		end
		$finish;
	end

endmodule





