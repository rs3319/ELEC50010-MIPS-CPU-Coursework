module ALU_32bit(
	
	input logic[5:0] ALU_control, opcode,
	input logic[4:0] shamt, // for shift
	input logic[15:0] immediate,
	input logic[31:0] rs_content, rt_content, //inputs
    input logic carry_in, //need this?
	
	output logic sig_branch, 
	output logic[31:0] ALU_result, //ALU outpu
    output logic carry_out, //need this?
    output logic zero
);	

	integer i; //for loop
	logic[31:0] temp; //sra command? 

	always_comb begin		
			
		// R-type instructions
		if(opcode == 6'h0) begin
			
			case(ALU_control)
				
				6'h21 : //addu
					ALU_result = rs_content + rt_content;
					
				6'h23 : //subu
					ALU_result = rs_content - rt_content;
					
				6'h24 : //and
					ALU_result = rs_content & rt_content;
					
				6'h25 : //or
					ALU_result = rs_content | rt_content;
					
				6'h03 : //sra
					begin
						temp = rt_content;
						for(i = 0; i < shamt; i = i + 1) begin
							temp = (temp[31],temp[31:1]); //add the lsb for msb
						end
					
					ALU_result = temp;
					end
					
				6'h02 : //srl
					ALU_result = (rt_content >> shamt);
			
				6'h00 : //sll
					ALU_result = (rt_content << shamt);
				
				6'h2b : //sltu
					begin
						if(rs_content < rt_content) begin
							ALU_result = 1;
						end 
                        else begin
							ALU_result = 0;
						end
					end
					
					end	
			endcase //case
			
		end // if		
		
		// I type instructions
		else begin
			
			signExtend = {{16{immediate[15]}}, immediate};
			zeroExtend = {{16{1'b0}}, immediate};
			
			case(opcode)
					
				6'h9 : // addiu
					ALU_result = rs_content + zeroExtend;
					
				6'b010010 : // andi
					ALU_result = rs_content & signExtend;
					
				6'h4 : // beq
					begin
						// if the result is zero, they are equal go branch
						ALU_result = rs_content - rt_content;
						if(ALU_result == 0) begin
							sig_branch = 1'b1;
						end
						else begin
							sig_branch = 1'b0;
						end
					end
				
				6'h5 : // bne
					begin
						// if the result is not zero, they are not equal go branch!
						ALU_result = rs_content - rt_content;
						if(ALU_result != 0) begin
							sig_branch = 1'b1;
							ALU_result = 1'b0;
						end
						else begin
							sig_branch = 1'b0;
						end
					end
				
				6'b010101 : // lui
					ALU_result = {immediate, {16{1'b0}};
				
				6'b010011 : // ori
					ALU_result = rs_content | zeroExtend;
				
				6'b001010 : // slti
					begin
						if($signed(rs_content) < $signed(signExtend)) begin
							ALU_result = 1;
						end else begin
							ALU_result = 0;
						end
					end
				
				6'b001011 : // sltiu
					begin
						if(rs_content < signExtend) begin
							ALU_result = 1;
						end else begin
							ALU_result = 0;
						end
					end
				
			endcase
		
		end
		
	end
	
	
	initial begin
		$monitor("opcode: %6b, Rs content: %32b, rt content: %32b, signExtendImm = %32b, result: %32b\n",
		opcode, rs_content, rt_content, signExtend, ALU_result);
	end
	
endmodule